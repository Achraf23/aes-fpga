----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07/14/2024 11:06:45 PM
-- Design Name: 
-- Module Name: top_TB - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity top_TB is
--  Port ( );
end top_TB;

architecture Behavioral of top_TB is
    component top is
        port (
            clk : in STD_LOGIC;
            out_bit : out STD_LOGIC
        );
    end component;
   
    signal sim_clk : std_logic := '0';
 
begin
    top_TB : top PORT MAP (
    clk=> sim_clk,
    out_bit => open
    );
    
    sim_clk <= not sim_clk after 5ns; 


end Behavioral;
